../../../rtl/vhdl/aes_top.vhdl