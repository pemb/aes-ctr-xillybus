../../../rtl/vhdl/aes_pkg.vhdl