../../../rtl/vhdl/colmix.vhdl