../../../rtl/vhdl/addkey.vhdl