../../../rtl/vhdl/mixcol.vhdl