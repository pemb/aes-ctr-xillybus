../../../rtl/vhdl/round.vhdl