../../../rtl/vhdl/subsh.vhdl