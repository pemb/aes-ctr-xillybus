../../../rtl/vhdl/keysched1.vhdl