../../../bench/vhdl/tb_aes.vhdl